module mux_2to1(i0, i1, sel, y);
    wire _0_;
    wire _1_;
    wire _2_;
    wire _3_;
    input i0;
    wire i0;
    input i1;
    wire i1;
    input sel;
    wire sel;
    output y;
    wire y;
    sky130_fd_sc_hd__mux2_1_4_ (
        .A0(_0_),
        .A1(_1_),
        .S(_2_),
        .X(_3_)
    );
    
    assign _0_ = i0;
    assign _1_ = i1;
    assign _2_ = sel;
    assign y = _3_;
endmodule
